module first_verilog_1 ();

wire    first_wire;
reg     first_reg;

assign  #10 first_wire = 1;

endmodule